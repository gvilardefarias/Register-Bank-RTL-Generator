`define ADDRESS_ADDR  12'h0
`define ADDRESS_STATUS  12'h4
