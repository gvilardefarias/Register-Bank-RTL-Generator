`define ADDRESS_ADDR  12'd0
`define ADDRESS_STATUS  12'd4
`define ADDRESS_MASK  12'd8
`define ADDRESS_DT_RCV  12'd12
`define ADDRESS_DT_TRA  12'd16
`define ADDRESS_DT_MX  12'd20
`define ADDRESS_WRITE_REG  12'd24
`define ADDRESS_READ_REG  12'd28
